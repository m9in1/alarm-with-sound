module sound_top(
	input clk,
	input rstn,
	input aud_en,
	output pwm

);



endmodule